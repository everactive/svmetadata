`include "uvm_pkg.sv"
`include "meta_pkg.sv"
