program svmetadata();
  initial uvm_pkg::run_test();
endprogram : svmetadata
